// Name: Leonard Paya, Rhiannon Garnier
// ID: 2200906, 2336462
// Due Date: 12/07/2025
// Class: EE 371


module pac_man_behavior_tb ();
    
    logic clk, reset;
    logic up, down, left, right;
    logic [9:0] curr_block;
    logic [9:0] next_block;

endmodule